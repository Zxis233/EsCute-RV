`include "include/defines.svh"
// [TODO] 实现乘法指令
// [HACK] 不阻塞EX级
// [HACK] 实现变长流水线
// [HACK] 实现华莱士树乘法器
