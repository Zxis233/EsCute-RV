`include "include/defines.svh"
// [TODO] 实现Zicsr扩展
